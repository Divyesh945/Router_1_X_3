/************************************************************************
  
Copyright 2019 - Maven Silicon Softech Pvt Ltd.  
  
www.maven-silicon.com 
  
All Rights Reserved. 
This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd. 
It is not to be shared with or used by any third parties who have not enrolled for our paid 
training courses or received any written authorization from Maven Silicon.
  
Filename:       ram_test_pkg.sv
  
Author Name:    Putta Satish

Support e-mail: For any queries, reach out to us on "techsupport_vm@maven-silicon.com" 

Version:	1.0

************************************************************************/
package router_test_pkg;


	//import uvm_pkg.sv
	import uvm_pkg::*;
	//include uvm_macros.sv
	`include "uvm_macros.svh"
	//`include "tb_defs.sv"
	`include "source_xtn.sv"
	`include "router_source_agent_config.sv"
	`include "router_destination_agent_config.sv"
	`include "router_env_config.sv"
	`include "router_source_driver.sv"
	`include "router_source_monitor.sv"
	`include "router_source_sequencer.sv"
	`include "router_source_agent.sv"
	`include "router_source_agt_top.sv"
	`include "router_source_seqs.sv"
	
	`include "destination_xtn.sv"
	`include "router_destination_monitor.sv"
	`include "router_destination_sequencer.sv"
	`include "router_destination_seqs.sv"
	`include "router_destination_driver.sv"
	`include "router_destination_agent.sv"
	`include "router_destination_agt_top.sv"
	
	`include "router_virtual_sequencer.sv"
	`include "router_virtual_seqs.sv"
	`include "router_sb.sv"
	
	`include "router_env.sv"
	
	
	`include "router_test.sv"
endpackage
